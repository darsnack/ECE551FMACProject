module multiplier(input CLK, input RESET,input [7:0] x, input [7:0] y, output [15:0] multOut);

