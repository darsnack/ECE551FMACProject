module adder12bit_behav(input [8:0] a, input [8:0] b, input cin, output cout, output [7:0] s);
