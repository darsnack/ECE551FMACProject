module multiplier(input [7:0] x, input [7:0] y, output [15:0] multOut);
	assign multOut = x*y;
endmodule
